netcdf example { // example of CDL notation
dimensions:
lon = 3 ;
lat = 8 ;
variables:
float rh(lon, lat) ;
rh:units = "percent" ;
rh:long_name = "Relative humidity" ;
// global attributes
:title = "Simple example, lacks some conventions" ;
data:
 rh =
 2, 3, 5, 7, 11, 13, 17, 19,
 23, 29, 31, 37, 41, 43, 47,
 53, 59, 61, 67, 71, 73, 79, 83, 89 ;
}
